0
49 58 61 215 19 g 38 47 43 55 60 54 46 37 30 21 13 29 26 20 12 9 5 3 6 1 0 2 7 10 14 18 22 31 35 39 52 63 67 69 71 70 65 61 c 37 3 25 3 30 1
4 7 7 5 10 g 56 48 64 c 32 2 44 1
9 4 3 7 0 g 24 50 33 41 58 62 59 51 c 16 2 40 1
1 0 2 0 0 g 27 32 c 20 1 27 1
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
9
