3
100 100 100 500 100 g 0 1 2 c 0 3 4 2
10 10 10 10 10 g 56 48 64 c 32 2 44 1
11 10 14 10 10 g 24 50 33 41 c 16 2 40 1
0 0 0 0 0 g 27 32 c 20 1 27 1
0 3 1 10 2 5 3 4 4 7 5 10 5 11 5 3 5 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
8
